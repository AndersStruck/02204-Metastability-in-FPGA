--------------------------------------------------------------------------------
--
-- Title    : hmw4.vhdl
-- Project  : Rounding
-- Author   : Jacob Jessen
-- Date     : Day/Month/YEAR
--------------------------------------------------------------------------------
--
-- Description
-- 
--------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
use IEEE.std_logic_signed.all;

hej

entity E is